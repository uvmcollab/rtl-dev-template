`ifndef VIF_IF_SV
`define VIF_IF_SV

interface vif_if(
    input logic clk_i
); 

  timeunit      1ns;
  timeprecision 1ps;
  
  localparam int Width = 8;

  logic rst_i;
  logic [Width-1:0] a_i;
  logic [Width-1:0] b_i;
  logic [Width-1:0] c_i;
  logic [Width-1:0] d_i;
  logic [Width-1:0] e_i;
  logic [Width-1:0] f_i;
  logic [Width-1:0] g_i;
  logic [Width-1:0] h_i;
  logic [Width-1:0] y_o;
  logic [2:0]sel_i;

  clocking cb @(posedge clk_i);
    default input #1ns output #1ns;
    output rst_i;
    output sel_i;
    output a_i;
    output b_i;
    output c_i;
    output d_i;
    output e_i;
    output f_i;
    output h_i;
    output g_i;
  endclocking : cb

endinterface : vif_if

`endif // VIF_IF_SV
