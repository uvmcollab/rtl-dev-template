// Design Code (DUT)
// FIFO

module fifo(
  input clk, rst, wr, rd, 
  input [7:0] din,
  output reg [7:0] dout,
  output reg empty, full);
  
  reg [3:0] wrop = 0,rdop = 0,cnt = 0;
  reg [7:0] mem [15:0];
  
  always@(posedge clk)
    begin
      if(rst== 1'b1)
         begin
           cnt <= 0;
           wrop <= 0;
           rdop= 0;
         end
      else if(wr && !full)
          begin
            if(cnt < 15) begin
              mem[wrop] <= din;
            wrop <= wrop + 1;
            cnt <= cnt + 1;
            end
          end
      else if (rd && !empty)
        begin
          if(cnt > 0) begin
            dout <= mem[rdop];
          rdop <= rdop + 1;
          cnt <= cnt - 1;
          end
        end 
      
      if(wrop == 15)
         wrop <= 0;
      if(rdop == 15)
         rdop <= 0;
    end
  
  assign empty = (cnt == 0) ? 1'b1 : 1'b0;
  assign full = (cnt == 15) ? 1'b1 : 1'b0;
  
endmodule